library verilog;
use verilog.vl_types.all;
entity majorita3_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end majorita3_vlg_check_tst;
