library verilog;
use verilog.vl_types.all;
entity KOM2_vlg_vec_tst is
end KOM2_vlg_vec_tst;
